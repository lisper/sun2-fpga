module ttl_am9513 (inout [15:0] D,
		   input  CD_n,
		   input  CS_n,
		   input  RD_n,
		   input  WR_n,
		   input  X1,
		   input  X2,
		   input  FOUT,
		   input  SRC1,
		   input  SRC2,
		   input  SRC3,
		   input  SRC4,
		   input  SRC5,
		   input  SRC6,
		   input  GAT1,
		   input  GAT2,
		   input  GAT3,
		   input  GAT4,
		   input  GAT5,
		   output OUT1,
		   output OUT2,
		   output OUT3,
		   output OUT4,
		   output OUT5);

   assign D = 16'bz;
   
endmodule

